library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity MyInstructionMemory is
       port (
       A  : in  STD_LOGIC_VECTOR(31 downto 0);
       RD : out STD_LOGIC_VECTOR(31 downto 0));
end MyInstructionMemory;

architecture Behavioral of MyInstructionMemory is
	type Memory is array (0 to 31) of STD_LOGIC_VECTOR(31 downto 0);
	signal IMem : Memory := (

      "10001100001000110000000000000010", --1 lw $t3, 2($t1) -- t3 = 1
      "10001100001001000000000000000010", --2 lw $t4, 2($t1) -- t4 = 1
      "00000000000000000000000000000000", --3 stall
      "00000000011001000010100000100000", --4 add $t5, $t3, $t4 -- 1 + 1
      "00000000000000000000000000000000", --5 stall
      "10101100001001010000000000000011", --6 sw $t5, 3($t1) -- 2 
      "10001100001001010000000000000011", --7 lw $t5, 3($t1) -- 2
      "00000000000000000000000000000000", --8 stall
      "00000000101001000011000000100000", --8 add $t6, $t5, $t4 -- 2 + 1
      "00000000000000000000000000000000", --9 stall
      "10101100001001100000000000000100", --10 sw $t6, 4($t1) -- 3 
      "10001100001001100000000000000100", --11 lw  $t6, 4($t1) -- 3
      "00000000000000000000000000000000", --12 stall
      "00000000101001100011100000100000", --13 add $t7, $t5, $t6 -- 2 + 3
      "00000000000000000000000000000000", --14 stall
      "10101100001001110000000000000101", --15 sw $t7, 5($t1) -- 5
      "10001100001001110000000000000101", --16 lw $t7, 5($t1) -- 5
      "00000000000000000000000000000000", --32 stall
      "00000000111001100100000000100000", --16 add $t8, $t7, $t6 -- 5 + 3
      "00000000000000000000000000000000", --17 stall
      "10101100001010000000000000000110", --18 sw $t8, 6($t1) -- 8
      "10001100001010000000000000000110", --19 lw $t8, 6($t1) -- 8
      "00000000000000000000000000000000", --32 stall
      "00000001000001110100100000100000", --20 add $t9, $t8, $t7 -- 8 + 5
      "00000000000000000000000000000000", --21 stall
      "10101100001010010000000000000111", --22 sw $t9, 7($t1) -- 13
      "10001100001010010000000000000111", --23 lw $t9, 7($t1) -- 13  
      "00000000000000000000000000000000", --28 stall
      "00000000000000000000000000000000", --29 stall
      "00000000000000000000000000000000", --30 stall
      "00000000000000000000000000000000", --31 stall
      "00000000000000000000000000000000" --32 stall
      );

begin

	process (A)
	begin
		RD <= IMem(TO_INTEGER(UNSIGNED(A)) / 4);
		
	end process;

end Behavioral;